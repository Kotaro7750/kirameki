package MulDivTypes;

import BasicTypes::*;
import OpTypes::*;

localparam MULDIV_PIPELINE_DEPTH = 5;

typedef logic [32:0] SignExtendedBasicData;
typedef logic [63:0] MulDivResult;

endpackage
