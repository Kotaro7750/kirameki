package ControllerTypes;
  typedef struct packed {
    logic stall;
    logic flush;
  } StageCtrl ;
endpackage
