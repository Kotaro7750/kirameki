//localparam CLOCKS_PER_SEC = 100000000;

//`define DEBUG

//`define BRANCH_M //条件分岐確定ステージ

`define NOT_USE_BTB //BTB使うのか
