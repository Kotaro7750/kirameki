//localparam CLOCKS_PER_SEC = 100000000;

`define DEBUG
//`define WITH_HC

//`define BRANCH_M //条件分岐確定ステージ

//`define BPRED_STATIC //静的分岐予測

//`define NOT_USE_BTB //BTB使うのか
